`include "uvm_macros.svh"
`include "top.sv"
